* SPICE3 file created from 5nand.ext - technology: scmos
.include TSMC_180nm.txt
.option scale=0.09u

M1000 a_54_n43# in4 a_28_n43# Gnd CMOSN w=10 l=2
+  ad=260 pd=72 as=240 ps=68
M1001 out in3 vdd w_n48_10# CMOSP w=10 l=2
+  ad=480 pd=196 as=470 ps=194
M1002 a_n29_n43# in1 gnd Gnd CMOSN w=10 l=2
+  ad=270 pd=74 as=90 ps=38
M1003 out in1 vdd w_n48_10# CMOSP w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1004 out in2 vdd w_n48_10# CMOSP w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1005 out in5 vdd w_n48_10# CMOSP w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1006 out in5 a_54_n43# Gnd CMOSN w=10 l=2
+  ad=100 pd=40 as=0 ps=0
M1007 a_0_n43# in2 a_n29_n43# Gnd CMOSN w=10 l=2
+  ad=260 pd=72 as=0 ps=0
M1008 out in4 vdd w_n48_10# CMOSP w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1009 a_28_n43# in3 a_0_n43# Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
C0 w_n48_10# Gnd 4.04fF

Vdd vdd gnd 2


V_in_a in1 gnd DC 2
V_in_b in2 gnd DC 2
V_in_c in3 gnd DC 2
V_in_d in4 gnd DC 2
V_in_e in5 gnd DC 2
.tran 1u 10000u




.control
run
set color0 = rgb:f/f/e
set color1 = black
plot v(out) v(in1)+3 v(in2)+5 v(in3)+7
.endc
.end