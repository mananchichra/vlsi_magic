magic
tech scmos
timestamp 1701035029
<< nwell >>
rect -14 2 22 23
<< ntransistor >>
rect 3 -13 5 -5
<< ptransistor >>
rect 3 8 5 16
<< ndiffusion >>
rect -8 -9 3 -5
rect -4 -13 3 -9
rect 5 -9 11 -5
rect 5 -13 15 -9
<< pdiffusion >>
rect -4 12 3 16
rect -8 8 3 12
rect 5 12 15 16
rect 5 8 11 12
<< ndcontact >>
rect -8 -13 -4 -9
rect 11 -9 15 -5
<< pdcontact >>
rect -8 12 -4 16
rect 11 8 15 12
<< polysilicon >>
rect 3 16 5 19
rect 3 -5 5 8
rect 3 -16 5 -13
<< polycontact >>
rect -1 -2 3 2
<< metal1 >>
rect -8 16 -5 23
rect -14 -2 -1 1
rect 12 -5 15 8
rect -8 -16 -5 -13
<< labels >>
rlabel metal1 -13 -1 -13 -1 3 in
rlabel metal1 14 0 14 0 1 out
rlabel metal1 -6 21 -6 21 5 vdd!
rlabel metal1 -7 -15 -7 -15 1 gnd!
<< end >>
