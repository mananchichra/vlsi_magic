magic
tech scmos
timestamp 1701502597
<< nwell >>
rect 4394 905 4430 926
rect 4459 918 4505 939
rect 4515 917 4551 938
rect 620 386 641 432
rect 1383 381 1404 427
rect 2159 384 2180 430
rect 619 340 640 376
rect 1382 335 1403 371
rect 2158 338 2179 374
<< ntransistor >>
rect 4475 902 4477 909
rect 4487 902 4489 909
rect 4532 902 4534 910
rect 4411 890 4413 898
rect 604 414 611 416
rect 2143 412 2150 414
rect 1367 409 1374 411
rect 604 402 611 404
rect 2143 400 2150 402
rect 1367 397 1374 399
rect 604 357 612 359
rect 2143 355 2151 357
rect 1367 352 1375 354
<< ptransistor >>
rect 4475 925 4477 932
rect 4487 925 4489 932
rect 4411 911 4413 919
rect 4532 923 4534 931
rect 627 414 634 416
rect 2166 412 2173 414
rect 1390 409 1397 411
rect 627 402 634 404
rect 2166 400 2173 402
rect 1390 397 1397 399
rect 625 357 633 359
rect 2164 355 2172 357
rect 1388 352 1396 354
<< ndiffusion >>
rect 4471 905 4475 909
rect 4467 902 4475 905
rect 4477 902 4487 909
rect 4489 905 4495 909
rect 4489 902 4499 905
rect 4521 906 4532 910
rect 4525 902 4532 906
rect 4534 906 4540 910
rect 4534 902 4544 906
rect 4400 894 4411 898
rect 4404 890 4411 894
rect 4413 894 4419 898
rect 4413 890 4423 894
rect 604 420 607 424
rect 604 416 611 420
rect 1367 415 1370 419
rect 604 404 611 414
rect 1367 411 1374 415
rect 2143 418 2146 422
rect 2143 414 2150 418
rect 604 396 611 402
rect 604 392 607 396
rect 1367 399 1374 409
rect 2143 402 2150 412
rect 1367 391 1374 397
rect 1367 387 1370 391
rect 2143 394 2150 400
rect 2143 390 2146 394
rect 608 366 612 370
rect 604 359 612 366
rect 1371 361 1375 365
rect 604 351 612 357
rect 604 347 608 351
rect 1367 354 1375 361
rect 2147 364 2151 368
rect 2143 357 2151 364
rect 1367 346 1375 352
rect 1367 342 1371 346
rect 2143 349 2151 355
rect 2143 345 2147 349
<< pdiffusion >>
rect 4470 928 4475 932
rect 4466 925 4475 928
rect 4477 930 4487 932
rect 4477 925 4480 930
rect 4485 925 4487 930
rect 4489 929 4498 932
rect 4489 925 4494 929
rect 4525 927 4532 931
rect 4404 915 4411 919
rect 4400 911 4411 915
rect 4413 915 4423 919
rect 4413 911 4419 915
rect 4521 923 4532 927
rect 4534 927 4544 931
rect 4534 923 4540 927
rect 627 421 630 425
rect 627 416 634 421
rect 1390 416 1393 420
rect 627 411 634 414
rect 1390 411 1397 416
rect 2166 419 2169 423
rect 2166 414 2173 419
rect 632 406 634 411
rect 627 404 634 406
rect 627 397 634 402
rect 1390 406 1397 409
rect 1395 401 1397 406
rect 2166 409 2173 412
rect 2171 404 2173 409
rect 2166 402 2173 404
rect 1390 399 1397 401
rect 631 393 634 397
rect 1390 392 1397 397
rect 1394 388 1397 392
rect 2166 395 2173 400
rect 2170 391 2173 395
rect 625 366 629 370
rect 625 359 633 366
rect 625 351 633 357
rect 1388 361 1392 365
rect 1388 354 1396 361
rect 2164 364 2168 368
rect 2164 357 2172 364
rect 629 347 633 351
rect 1388 346 1396 352
rect 1392 342 1396 346
rect 2164 349 2172 355
rect 2168 345 2172 349
<< ndcontact >>
rect 4467 905 4471 909
rect 4495 905 4499 909
rect 4521 902 4525 906
rect 4540 906 4544 910
rect 4400 890 4404 894
rect 4419 894 4423 898
rect 607 420 611 424
rect 1370 415 1374 419
rect 2146 418 2150 422
rect 607 392 611 396
rect 1370 387 1374 391
rect 2146 390 2150 394
rect 604 366 608 370
rect 1367 361 1371 365
rect 608 347 612 351
rect 2143 364 2147 368
rect 1371 342 1375 346
rect 2147 345 2151 349
<< pdcontact >>
rect 4466 928 4470 932
rect 4494 925 4498 929
rect 4521 927 4525 931
rect 4400 915 4404 919
rect 4419 911 4423 915
rect 4540 923 4544 927
rect 630 421 634 425
rect 1393 416 1397 420
rect 2169 419 2173 423
rect 627 393 631 397
rect 1390 388 1394 392
rect 2166 391 2170 395
rect 629 366 633 370
rect 1392 361 1396 365
rect 2168 364 2172 368
rect 625 347 629 351
rect 1388 342 1392 346
rect 2164 345 2168 349
<< polysilicon >>
rect 4475 932 4477 935
rect 4487 932 4489 935
rect 4532 931 4534 934
rect 4411 919 4413 922
rect 4411 898 4413 911
rect 4475 909 4477 925
rect 4487 909 4489 925
rect 4532 910 4534 923
rect 4475 899 4477 902
rect 4487 899 4489 902
rect 4532 899 4534 902
rect 4411 887 4413 890
rect 601 414 604 416
rect 611 414 627 416
rect 634 414 637 416
rect 2140 412 2143 414
rect 2150 412 2166 414
rect 2173 412 2176 414
rect 1364 409 1367 411
rect 1374 409 1390 411
rect 1397 409 1400 411
rect 601 402 604 404
rect 611 402 627 404
rect 634 402 637 404
rect 2140 400 2143 402
rect 2150 400 2166 402
rect 2173 400 2176 402
rect 1364 397 1367 399
rect 1374 397 1390 399
rect 1397 397 1400 399
rect 601 357 604 359
rect 612 357 625 359
rect 633 357 636 359
rect 2140 355 2143 357
rect 2151 355 2164 357
rect 2172 355 2175 357
rect 1364 352 1367 354
rect 1375 352 1388 354
rect 1396 352 1399 354
<< polycontact >>
rect 4471 920 4475 924
rect 4407 901 4411 905
rect 4483 914 4487 918
rect 4528 913 4532 917
rect 622 416 626 420
rect 1385 411 1389 415
rect 2161 414 2165 418
rect 616 404 620 408
rect 1379 399 1383 403
rect 2155 402 2159 406
rect 615 359 619 363
rect 1378 354 1382 358
rect 2154 357 2158 361
<< metal1 >>
rect 3574 982 4629 985
rect 3596 773 3599 982
rect 4383 951 4433 956
rect 4439 951 4444 954
rect 4383 828 4388 951
rect 4400 919 4403 925
rect 4441 924 4444 951
rect 4469 936 4498 939
rect 4469 932 4472 936
rect 4470 928 4472 932
rect 4481 930 4484 932
rect 4495 929 4498 936
rect 4521 931 4524 934
rect 4441 921 4471 924
rect 4495 921 4498 925
rect 4495 918 4514 921
rect 4399 901 4407 904
rect 4420 903 4423 911
rect 4435 914 4483 917
rect 4435 903 4438 914
rect 4495 909 4498 918
rect 4511 916 4514 918
rect 4541 917 4544 923
rect 4511 913 4528 916
rect 4541 914 4547 917
rect 4541 910 4544 914
rect 4420 900 4438 903
rect 4544 906 4545 909
rect 4420 898 4423 900
rect 4467 899 4470 905
rect 4521 899 4524 902
rect 4467 896 4524 899
rect 4398 890 4400 891
rect 4511 891 4514 896
rect 4404 890 4514 891
rect 4398 888 4514 890
rect 4400 887 4403 888
rect 4511 829 4514 888
rect 4542 886 4545 906
rect 4626 886 4629 982
rect 4542 883 4654 886
rect 4542 877 4545 883
rect 4383 823 4389 828
rect 4511 826 4651 829
rect 4412 816 4438 819
rect 4392 805 4395 807
rect 3367 772 3599 773
rect 4369 802 4395 805
rect 3367 771 3618 772
rect 3367 769 3619 771
rect 3367 768 3612 769
rect 3367 569 3370 768
rect 3616 764 3619 766
rect 3590 761 3619 764
rect 3708 762 3715 765
rect 3590 709 3593 761
rect 4369 756 4372 802
rect 4435 789 4438 816
rect 4435 786 4453 789
rect 4429 779 4459 782
rect 4429 768 4432 779
rect 4537 772 4539 774
rect 4414 765 4432 768
rect 4505 756 4508 764
rect 4369 753 4508 756
rect 3525 706 3593 709
rect 3495 675 3498 691
rect 3672 675 3675 747
rect 3495 672 3689 675
rect 3367 567 3574 569
rect 3367 566 3582 567
rect 23 495 652 501
rect 23 427 29 495
rect 71 474 73 475
rect 646 451 652 495
rect 3523 476 3526 566
rect 3571 564 3582 566
rect 3573 557 3581 560
rect 3666 557 3677 560
rect 3523 473 3541 476
rect 646 445 2198 451
rect 646 443 660 445
rect 616 433 619 434
rect 571 430 619 433
rect 4 421 50 427
rect 4 392 10 421
rect -130 386 10 392
rect -130 59 -124 386
rect 64 360 68 384
rect -103 356 68 360
rect -103 170 -99 356
rect 571 325 574 430
rect 598 421 607 424
rect 598 385 601 421
rect 616 408 619 430
rect 623 420 626 434
rect 634 421 641 422
rect 630 419 641 421
rect 632 407 634 410
rect 611 393 627 396
rect 638 396 641 419
rect 631 393 641 396
rect 583 381 601 385
rect 583 334 587 381
rect 598 370 601 381
rect 620 380 623 393
rect 615 377 623 380
rect 598 367 604 370
rect 615 363 618 377
rect 633 367 636 370
rect 612 347 625 350
rect 616 338 619 347
rect 654 334 660 443
rect 1379 426 1382 429
rect 583 330 660 334
rect 1343 423 1383 426
rect 571 322 672 325
rect 669 177 672 322
rect 1343 280 1346 423
rect 1361 416 1370 419
rect 1361 373 1364 416
rect 1379 403 1382 423
rect 1386 415 1389 428
rect 1397 416 1404 417
rect 1393 414 1404 416
rect 1395 402 1397 405
rect 1374 388 1390 391
rect 1401 391 1404 414
rect 1394 388 1404 391
rect 1383 375 1386 388
rect 1354 369 1364 373
rect 1354 326 1358 369
rect 1361 365 1364 369
rect 1378 372 1386 375
rect 1361 362 1367 365
rect 1378 358 1381 372
rect 1396 362 1399 365
rect 1375 342 1388 345
rect 1379 336 1382 342
rect 1437 326 1443 445
rect 2110 431 2158 434
rect 1354 320 1443 326
rect 2110 322 2113 431
rect 2137 419 2146 422
rect 2137 385 2140 419
rect 2155 406 2158 431
rect 2162 418 2165 431
rect 2173 419 2180 420
rect 2169 417 2180 419
rect 2171 405 2173 408
rect 2150 391 2166 394
rect 2177 394 2180 417
rect 2170 391 2180 394
rect 2120 379 2142 385
rect 2120 334 2126 379
rect 2137 368 2140 379
rect 2159 378 2162 391
rect 2154 375 2162 378
rect 2137 365 2143 368
rect 2154 361 2157 375
rect 2172 365 2175 368
rect 2151 345 2164 348
rect 2155 337 2158 345
rect 2192 334 2198 445
rect 3538 338 3541 473
rect 3573 408 3576 557
rect 3627 536 3630 542
rect 3686 536 3689 672
rect 3627 533 3689 536
rect 4505 534 4508 753
rect 4536 707 4539 772
rect 4536 704 4545 707
rect 4536 657 4539 704
rect 4633 697 4642 700
rect 4648 682 4651 826
rect 4611 679 4651 682
rect 4536 654 4546 657
rect 4536 605 4539 654
rect 4632 647 4640 650
rect 4648 632 4651 679
rect 4609 629 4651 632
rect 4536 602 4543 605
rect 4632 595 4639 598
rect 4648 580 4651 629
rect 3686 442 3689 533
rect 4555 532 4558 580
rect 4606 577 4651 580
rect 3686 439 3718 442
rect 3715 428 3718 439
rect 3715 425 3748 428
rect 3573 405 3669 408
rect 3666 372 3669 405
rect 3661 369 3669 372
rect 3630 351 3792 354
rect 2120 328 2198 334
rect 3434 335 3593 338
rect 2110 319 2215 322
rect 1343 277 1401 280
rect 1398 238 1401 277
rect 1398 235 1456 238
rect 1453 174 1456 235
rect 2212 177 2215 319
rect 3024 196 3026 197
rect 2983 193 3027 196
rect 3115 194 3124 197
rect 3434 195 3437 335
rect 3590 291 3593 335
rect 3590 288 3647 291
rect 3644 250 3647 288
rect 3644 247 3655 250
rect 3637 241 3655 244
rect 3741 241 3751 244
rect 3637 231 3640 241
rect 3560 228 3640 231
rect 3701 213 3704 226
rect 3835 213 3838 266
rect 3531 210 3838 213
rect 3701 209 3704 210
rect 2983 174 2986 193
rect 3434 192 3608 195
rect -103 166 -61 170
rect -65 84 -61 166
rect 3605 163 3608 192
rect 3592 160 3608 163
rect 3592 107 3595 160
rect 3003 102 3040 105
rect 3122 102 3129 105
rect 3592 104 3614 107
rect 3003 96 3007 102
rect 3600 97 3607 100
rect 3696 97 3704 100
rect 2988 92 3007 96
rect 3600 88 3603 97
rect -65 80 -48 84
rect 3567 85 3603 88
rect 3533 67 3616 70
rect 3651 70 3654 82
rect 4046 70 4049 76
rect 3622 67 4049 70
rect -130 53 -46 59
<< m2contact >>
rect 4433 951 4439 957
rect 4400 925 4405 930
rect 4520 934 4525 939
rect 4394 901 4399 906
rect 4392 841 4397 846
rect 4386 818 4391 823
rect 3433 713 3438 718
rect 4394 790 4399 795
rect 4388 766 4393 771
rect 3435 704 3440 709
rect 63 473 68 478
rect 73 472 78 477
rect 623 434 628 439
rect 636 366 641 371
rect 1386 428 1391 433
rect 1399 361 1404 366
rect 2162 431 2167 436
rect 2175 364 2180 369
rect 4479 614 4484 619
rect 4441 590 4446 595
rect 4493 562 4498 567
rect 4545 696 4550 701
rect 4542 645 4547 650
rect 4542 594 4547 599
rect 3569 376 3574 381
rect 3568 367 3573 372
rect 3020 200 3025 205
rect 3468 235 3473 240
rect 3467 226 3472 231
rect 3029 108 3034 113
rect 3475 92 3480 97
rect 3475 83 3480 88
<< pdm12contact >>
rect 4480 925 4485 930
rect 627 406 632 411
rect 1390 401 1395 406
rect 2166 404 2171 409
<< metal2 >>
rect 4080 953 4433 956
rect 4080 952 4359 953
rect 4080 878 4084 952
rect 4466 946 4469 952
rect 4465 943 4469 946
rect 4465 937 4468 943
rect 4511 942 4587 945
rect 4511 937 4514 942
rect 4520 939 4525 942
rect 4449 934 4520 937
rect 4412 929 4415 930
rect 4449 929 4452 934
rect 4481 930 4484 934
rect 4405 926 4452 929
rect 63 874 4084 878
rect 4102 901 4394 904
rect 63 478 67 874
rect 4102 863 4105 901
rect 77 860 4105 863
rect 77 481 80 860
rect 3487 736 3609 737
rect 3670 736 3673 785
rect 4339 769 4342 901
rect 4397 843 4463 846
rect 4385 818 4386 821
rect 4406 794 4409 843
rect 4460 811 4463 843
rect 4459 808 4463 811
rect 4580 810 4583 942
rect 4505 807 4591 810
rect 4505 799 4508 807
rect 4514 804 4519 807
rect 4399 791 4409 794
rect 4338 766 4388 769
rect 3487 734 3673 736
rect 3487 726 3490 734
rect 3498 730 3504 734
rect 3606 733 3673 734
rect 4588 736 4591 807
rect 4588 733 4596 736
rect 3400 714 3433 718
rect 3400 656 3404 714
rect 3432 713 3433 714
rect 3422 706 3435 709
rect 3422 670 3425 706
rect 3440 706 3443 709
rect 3606 693 3609 733
rect 4593 720 4596 733
rect 4592 718 4596 720
rect 4441 696 4545 701
rect 3606 690 3732 693
rect 3729 673 3732 690
rect 3729 670 3844 673
rect 3422 661 3426 664
rect 3400 644 3404 650
rect 3627 596 3684 600
rect 3627 578 3631 596
rect 3680 580 3684 596
rect 4441 595 4446 696
rect 4484 650 4543 651
rect 4484 646 4542 650
rect 4484 614 4489 646
rect 4592 620 4595 718
rect 4494 594 4542 599
rect 3680 576 3843 580
rect 4494 567 4499 594
rect 4591 571 4595 620
rect 4591 567 4603 571
rect 75 477 628 481
rect 78 475 80 477
rect 624 440 628 477
rect 624 439 3031 440
rect 628 436 3031 439
rect 1381 433 2162 436
rect 2167 433 3031 436
rect 84 421 154 424
rect 151 313 154 421
rect 636 423 645 426
rect 636 410 639 423
rect 2175 421 2184 424
rect 632 407 639 410
rect 636 383 639 407
rect 1399 418 1408 421
rect 1399 405 1402 418
rect 1395 402 1402 405
rect 2175 408 2178 421
rect 2171 405 2178 408
rect 636 380 691 383
rect 636 371 639 380
rect 688 312 691 380
rect 1399 378 1402 402
rect 2175 380 2178 405
rect 1399 375 1423 378
rect 1399 366 1402 375
rect 1420 312 1423 375
rect 2175 377 2193 380
rect 2175 369 2178 377
rect 2190 311 2193 377
rect 3021 258 3028 433
rect 3553 371 3557 463
rect 3597 428 3601 514
rect 4599 498 4603 567
rect 4513 494 4603 498
rect 3562 424 3601 428
rect 3562 385 3566 424
rect 3562 376 3569 385
rect 3553 367 3568 371
rect 3624 341 3627 393
rect 3703 341 3706 342
rect 3624 338 3878 341
rect 3448 328 3497 332
rect 3001 251 3156 258
rect 3001 206 3008 251
rect 3001 205 3022 206
rect 3001 200 3020 205
rect 3001 199 3022 200
rect 3072 193 3075 217
rect 3049 190 3075 193
rect 3049 163 3052 190
rect 3040 160 3052 163
rect 2868 135 2898 138
rect 3040 135 3043 160
rect 2866 132 2869 135
rect 2894 132 3043 135
rect 3040 131 3043 132
rect 3034 108 3035 112
rect 2710 60 2835 63
rect 2832 32 2835 60
rect 3031 58 3035 108
rect 3149 58 3156 251
rect 3448 231 3452 328
rect 3493 326 3497 328
rect 3526 317 3530 320
rect 3527 298 3530 317
rect 3499 295 3530 298
rect 3499 274 3502 295
rect 3624 276 3627 338
rect 3465 271 3502 274
rect 3520 273 3627 276
rect 3465 235 3468 271
rect 3520 248 3523 273
rect 3473 235 3478 238
rect 3448 227 3467 231
rect 3624 208 3627 273
rect 3579 205 3627 208
rect 3463 183 3464 185
rect 3458 182 3464 183
rect 3458 177 3465 182
rect 3435 85 3439 157
rect 3458 99 3464 177
rect 3579 141 3582 205
rect 3703 194 3706 338
rect 3528 138 3582 141
rect 3658 191 3706 194
rect 3658 140 3661 191
rect 3528 104 3531 138
rect 3657 137 3748 140
rect 3658 117 3661 137
rect 3458 97 3484 99
rect 3458 93 3475 97
rect 3480 93 3484 97
rect 3468 85 3475 88
rect 3435 83 3475 85
rect 3435 81 3476 83
rect 3030 51 3156 58
rect 3745 32 3748 137
rect 2832 29 3748 32
<< m3contact >>
rect 3421 664 3427 670
rect 3400 650 3406 656
rect 3597 514 3603 520
rect 3552 463 3558 469
rect 3497 326 3503 332
rect 3526 320 3532 326
rect 3457 183 3463 189
rect 3433 157 3439 163
<< m123contact >>
rect 4094 663 4099 668
rect 4091 634 4096 639
rect 4092 515 4097 520
rect 84 323 89 328
rect 102 324 107 329
rect 718 322 723 327
rect 739 325 744 330
rect 1461 323 1466 328
rect 1480 326 1485 331
rect 2230 326 2235 331
rect 2252 327 2257 332
rect 4087 463 4092 468
rect 3073 175 3078 180
rect 3084 83 3089 88
rect 4092 320 4097 325
rect 4090 306 4095 311
rect 4089 160 4094 165
rect 4080 153 4085 158
rect 3616 67 3622 72
<< metal3 >>
rect 184 665 3421 668
rect 184 363 187 665
rect 3427 666 3556 668
rect 4091 666 4094 668
rect 3427 665 4094 666
rect 3540 663 4094 665
rect 3540 662 3563 663
rect 81 360 187 363
rect 200 650 3400 655
rect 3406 650 3500 655
rect 81 332 84 360
rect 102 334 107 337
rect 200 334 205 650
rect 3495 641 3500 650
rect 3495 638 3541 641
rect 4088 638 4091 639
rect 3495 636 4091 638
rect 3495 629 3500 636
rect 3533 635 4091 636
rect 4088 634 4091 635
rect 81 329 89 332
rect 84 328 89 329
rect 102 329 205 334
rect 721 609 3547 614
rect 721 328 726 609
rect 741 587 2017 590
rect 741 584 3497 587
rect 741 580 2017 584
rect 741 330 751 580
rect 716 327 726 328
rect 716 323 718 327
rect 723 323 726 327
rect 744 325 751 330
rect 1462 533 3424 536
rect 1462 328 1465 533
rect 1483 489 3383 492
rect 1483 331 1486 489
rect 1485 327 1486 331
rect 2230 447 3273 452
rect 2230 331 2235 447
rect 2254 421 3221 425
rect 2254 332 2258 421
rect 2257 330 2258 332
rect 3217 299 3221 421
rect 3268 329 3273 447
rect 3380 406 3383 489
rect 3421 430 3424 533
rect 3494 468 3497 584
rect 3542 520 3547 609
rect 3537 515 3597 520
rect 3603 515 4092 520
rect 3494 465 3552 468
rect 3558 465 4087 468
rect 4084 464 4087 465
rect 3421 427 3529 430
rect 3380 403 3501 406
rect 3498 332 3501 403
rect 3268 324 3408 329
rect 3526 326 3529 427
rect 3217 295 3349 299
rect 3074 159 3077 175
rect 3345 162 3349 295
rect 3403 188 3408 324
rect 3498 311 3501 326
rect 3532 320 4092 323
rect 3498 308 4090 311
rect 4087 307 4090 308
rect 3403 183 3457 188
rect 3463 183 4090 188
rect 4086 172 4090 183
rect 4086 167 4092 172
rect 4089 165 4092 167
rect 3074 156 3087 159
rect 3345 158 3433 162
rect 3439 160 4081 162
rect 3439 158 4083 160
rect 4078 157 4080 158
rect 3084 88 3087 156
rect 3085 68 3089 83
rect 2937 64 3089 68
rect 2950 47 2954 64
rect 3617 47 3621 67
rect 2950 43 3621 47
use and2  and2_12
timestamp 1701462821
transform 1 0 3654 0 1 225
box -2 -2 92 45
use and2  and2_11
timestamp 1701462821
transform 1 0 3609 0 1 81
box -2 -2 92 45
use and2  and2_9
timestamp 1701462821
transform 1 0 3573 0 1 353
box -2 -2 92 45
use and2  and2_8
timestamp 1701462821
transform 1 0 3472 0 1 212
box -2 -2 92 45
use and2  and2_7
timestamp 1701462821
transform 1 0 3479 0 1 69
box -2 -2 92 45
use full_adder  full_adder_0
timestamp 1701449886
transform 1 0 23 0 1 5
box -105 13 2966 329
use and2  and2_0
timestamp 1701462821
transform 0 1 48 -1 0 472
box -2 -2 92 45
use and2  and2_2
timestamp 1701462821
transform 1 0 3027 0 1 178
box -2 -2 92 45
use and2  and2_3
timestamp 1701462821
transform 1 0 3034 0 1 86
box -2 -2 92 45
use and2  and2_14
timestamp 1701462821
transform 1 0 3579 0 1 541
box -2 -2 92 45
use and2  and2_13
timestamp 1701462821
transform 1 0 3620 0 1 746
box -2 -2 92 45
use and2  and2_10
timestamp 1701462821
transform 1 0 3437 0 1 690
box -2 -2 92 45
use not  not_1
timestamp 1701035029
transform 1 0 4402 0 1 768
box -14 -16 22 23
use and2  and2_1
timestamp 1701462821
transform 1 0 4544 0 1 631
box -2 -2 92 45
use and2  and2_4
timestamp 1701462821
transform 1 0 4544 0 1 579
box -2 -2 92 45
use and2  and2_5
timestamp 1701462821
transform 1 0 4546 0 1 681
box -2 -2 92 45
use and2  and2_6
timestamp 1701462821
transform 1 0 4453 0 1 763
box -2 -2 92 45
use not  not_0
timestamp 1701035029
transform 1 0 4400 0 1 820
box -14 -16 22 23
use comparator2  comparator2_0
timestamp 1701288896
transform 1 0 4221 0 1 476
box -521 -411 337 289
<< labels >>
rlabel metal1 4637 596 4637 596 1 b_gr
rlabel metal1 4638 648 4638 648 1 a_gr
rlabel metal1 4636 697 4642 700 1 equal
rlabel metal2 4105 953 4105 953 1 select0
rlabel metal2 4113 903 4113 903 1 select1
rlabel metal3 3253 666 3253 666 1 b0
rlabel metal3 3279 651 3279 651 1 a0
rlabel metal3 3271 611 3271 611 1 b1
rlabel metal3 3296 586 3296 586 1 a1
rlabel metal3 3302 534 3302 534 1 b2
rlabel metal3 3343 490 3343 490 1 a2
rlabel metal3 3304 326 3304 326 1 b3
rlabel metal3 3350 161 3350 161 1 a3
rlabel metal1 -125 55 -125 55 3 gnd!
rlabel metal2 2834 30 2834 31 1 vdd!
rlabel metal1 617 339 617 340 1 s0
rlabel metal1 1381 337 1381 338 1 s1
rlabel metal1 2156 339 2156 340 1 s2
rlabel metal1 3122 196 3122 197 1 s3
rlabel metal1 3128 103 3128 103 1 c_out
rlabel metal1 3703 98 3703 98 1 ab3
rlabel metal1 3750 242 3750 242 1 ab2
rlabel metal1 3675 558 3675 558 1 ab1
rlabel metal1 3713 763 3713 763 1 ab0
<< end >>
