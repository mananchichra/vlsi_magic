magic
tech scmos
timestamp 1701449886
<< metal1 >>
rect -105 306 -38 311
rect 62 299 66 324
rect -105 295 66 299
rect -105 245 -101 295
rect 80 292 84 325
rect -83 288 84 292
rect -83 265 -79 288
rect -86 261 -26 265
rect -105 241 -70 245
rect -74 176 -70 241
rect -86 172 -31 176
rect 659 172 663 175
rect 696 173 700 325
rect 716 278 719 325
rect 716 275 763 278
rect 760 258 763 275
rect 1439 272 1443 328
rect 1457 286 1461 327
rect 1457 282 1487 286
rect 1439 268 1472 272
rect 1468 176 1472 268
rect 1483 265 1487 282
rect 2207 273 2211 327
rect 2230 318 2235 329
rect 2230 279 2234 318
rect 2230 275 2258 279
rect 2207 269 2226 273
rect 1483 261 1511 265
rect -78 171 -74 172
rect 696 169 753 173
rect 1468 172 1504 176
rect 2200 172 2203 175
rect 2222 173 2226 269
rect 2254 262 2258 275
rect 2254 258 2269 262
rect 1445 169 1452 172
rect -44 165 -39 169
rect -86 164 -39 165
rect -34 164 -31 165
rect -86 161 -41 164
rect 1468 135 1472 172
rect 2221 169 2265 173
rect 2958 169 2966 172
rect 2221 122 2225 169
rect 658 90 756 94
rect -78 75 -37 79
rect 752 72 756 90
rect 1444 87 1511 91
rect 2199 90 2282 94
rect 1507 75 1511 87
rect 2278 72 2282 90
rect 2962 87 2966 91
rect -78 48 -34 54
rect 70 48 74 54
<< metal2 >>
rect 475 305 2356 310
rect 484 304 840 305
rect 1265 302 1585 305
<< m123contact >>
rect -39 164 -34 169
rect 745 161 750 166
rect 1500 164 1505 169
rect 2258 161 2263 166
<< metal3 >>
rect -39 298 2240 301
rect -39 169 -36 298
rect 738 164 741 298
rect 1484 168 1487 298
rect 738 161 745 164
rect 1484 165 1500 168
rect 2237 163 2240 298
rect 2237 161 2258 163
rect 2237 160 2261 161
rect 1261 20 1846 24
rect 468 16 1088 20
rect 2014 16 2607 20
use half_adder  half_adder_3
timestamp 1701446779
transform 1 0 2286 0 1 91
box -27 -78 676 217
use half_adder  half_adder_2
timestamp 1701446779
transform 1 0 1527 0 1 94
box -27 -78 676 217
use half_adder  half_adder_1
timestamp 1701446779
transform 1 0 772 0 1 91
box -27 -78 676 217
use half_adder  half_adder_0
timestamp 1701446779
transform 1 0 -14 0 1 94
box -27 -78 676 217
<< labels >>
rlabel metal1 65 320 65 323 5 b0
rlabel metal1 82 321 82 321 1 a0
rlabel metal1 697 320 697 320 1 b1
rlabel metal1 718 321 718 321 1 a1
rlabel metal1 1459 321 1459 321 1 a2
rlabel metal1 1441 323 1441 323 1 b2
rlabel metal1 2209 322 2209 322 1 b3
rlabel metal1 2233 323 2233 323 1 a3
rlabel metal1 2963 170 2963 170 7 s3
rlabel metal1 -82 163 -82 163 1 m
rlabel metal1 -76 77 -76 77 1 cin
rlabel metal1 -102 308 -102 308 3 vdd!
rlabel metal1 -74 50 -74 50 1 gnd!
rlabel metal1 2964 89 2964 89 7 c_out
rlabel metal1 2202 173 2202 173 1 s2
rlabel metal1 1448 170 1448 170 1 s1
rlabel metal1 661 174 661 174 1 s0
<< end >>
