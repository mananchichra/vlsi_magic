magic
tech scmos
timestamp 1701275880
<< nwell >>
rect 2 -52 80 -32
<< ntransistor >>
rect 13 -81 15 -75
rect 29 -81 31 -75
rect 47 -81 49 -75
rect 65 -81 67 -75
<< ptransistor >>
rect 13 -45 15 -38
rect 29 -45 31 -38
rect 47 -45 49 -38
rect 65 -45 67 -38
<< ndiffusion >>
rect 8 -77 13 -75
rect 12 -81 13 -77
rect 15 -81 29 -75
rect 31 -81 47 -75
rect 49 -81 65 -75
rect 67 -79 68 -75
rect 67 -81 72 -79
<< pdiffusion >>
rect 12 -42 13 -38
rect 8 -45 13 -42
rect 15 -41 20 -38
rect 15 -45 16 -41
rect 28 -42 29 -38
rect 24 -45 29 -42
rect 31 -41 37 -38
rect 31 -45 33 -41
rect 41 -42 42 -38
rect 46 -42 47 -38
rect 41 -45 47 -42
rect 49 -41 54 -38
rect 49 -45 50 -41
rect 59 -42 60 -38
rect 64 -42 65 -38
rect 59 -45 65 -42
rect 67 -41 72 -38
rect 67 -45 68 -41
<< ndcontact >>
rect 8 -81 12 -77
rect 68 -79 72 -75
<< pdcontact >>
rect 8 -42 12 -38
rect 16 -45 20 -41
rect 24 -42 28 -38
rect 33 -45 37 -41
rect 42 -42 46 -38
rect 50 -45 54 -41
rect 60 -42 64 -38
rect 68 -45 72 -41
<< polysilicon >>
rect 13 -38 15 -35
rect 29 -38 31 -35
rect 47 -38 49 -35
rect 65 -38 67 -35
rect 13 -75 15 -45
rect 29 -75 31 -45
rect 47 -75 49 -45
rect 65 -75 67 -45
rect 13 -84 15 -81
rect 29 -84 31 -81
rect 47 -84 49 -81
rect 65 -84 67 -81
<< polycontact >>
rect 9 -51 13 -47
rect 25 -58 29 -54
rect 43 -66 47 -62
rect 61 -73 65 -69
<< metal1 >>
rect 2 -32 63 -29
rect 8 -38 11 -32
rect 24 -38 27 -32
rect 42 -38 45 -32
rect 60 -38 63 -32
rect 2 -51 9 -48
rect 17 -48 72 -45
rect 2 -57 25 -54
rect 2 -65 43 -62
rect 2 -72 61 -69
rect 69 -75 72 -48
rect 8 -84 11 -81
<< labels >>
rlabel metal1 3 -31 3 -31 4 vdd!
rlabel metal1 3 -50 3 -50 3 in1
rlabel metal1 10 -83 10 -83 1 gnd!
rlabel metal1 71 -60 71 -60 1 out
rlabel metal1 4 -55 4 -55 3 in2
rlabel metal1 3 -63 3 -63 3 in3
rlabel metal1 3 -71 3 -71 3 in4
<< end >>
