magic
tech scmos
timestamp 1701462821
<< metal1 >>
rect -2 23 1 26
rect 49 20 55 23
rect -2 16 1 19
rect 52 18 55 20
rect 52 15 58 18
rect 85 16 88 19
rect 8 -2 65 1
<< m2contact >>
rect 61 36 66 41
<< metal2 >>
rect 6 41 9 45
rect 25 36 61 39
use not  not_0
timestamp 1701035029
transform 1 0 70 0 1 17
box -14 -16 22 23
use 2nand  2nand_0
timestamp 1700774385
transform 1 0 39 0 1 3
box -39 -3 10 38
<< labels >>
rlabel metal1 -1 24 -1 24 3 in1
rlabel metal1 -1 17 -1 17 3 in2
rlabel metal1 87 17 87 17 7 out
rlabel metal2 7 44 7 44 5 vdd!
rlabel metal1 64 -1 64 -1 1 gnd!
<< end >>
