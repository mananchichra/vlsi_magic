magic
tech scmos
timestamp 1701034208
<< nwell >>
rect -48 10 101 37
<< ntransistor >>
rect -31 -43 -29 -33
rect -2 -43 0 -33
rect 26 -43 28 -33
rect 52 -43 54 -33
rect 80 -43 82 -33
<< ptransistor >>
rect -31 18 -29 28
rect -2 18 0 28
rect 26 18 28 28
rect 52 18 54 28
rect 80 18 82 28
<< ndiffusion >>
rect -40 -39 -31 -33
rect -36 -43 -31 -39
rect -29 -43 -2 -33
rect 0 -43 26 -33
rect 28 -43 52 -33
rect 54 -43 80 -33
rect 82 -37 88 -33
rect 82 -43 92 -37
<< pdiffusion >>
rect -36 24 -31 28
rect -40 18 -31 24
rect -29 22 -19 28
rect -29 18 -23 22
rect -8 24 -2 28
rect -12 18 -2 24
rect 0 22 9 28
rect 0 18 5 22
rect 20 24 26 28
rect 16 18 26 24
rect 28 22 37 28
rect 28 18 33 22
rect 47 24 52 28
rect 43 18 52 24
rect 54 22 64 28
rect 54 18 60 22
rect 75 24 80 28
rect 71 18 80 24
rect 82 22 92 28
rect 82 18 88 22
<< ndcontact >>
rect -40 -43 -36 -39
rect 88 -37 92 -33
<< pdcontact >>
rect -40 24 -36 28
rect -23 18 -19 22
rect -12 24 -8 28
rect 5 18 9 22
rect 16 24 20 28
rect 33 18 37 22
rect 43 24 47 28
rect 60 18 64 22
rect 71 24 75 28
rect 88 18 92 22
<< polysilicon >>
rect -31 28 -29 31
rect -2 28 0 31
rect 26 28 28 31
rect 52 28 54 31
rect 80 28 82 31
rect -31 -33 -29 18
rect -2 -33 0 18
rect 26 -33 28 18
rect 52 -33 54 18
rect 80 -33 82 18
rect -31 -46 -29 -43
rect -2 -46 0 -43
rect 26 -46 28 -43
rect 52 -46 54 -43
rect 80 -46 82 -43
<< polycontact >>
rect -35 7 -31 11
rect -6 -2 -2 2
rect 22 -10 26 -6
rect 48 -19 52 -15
rect 76 -28 80 -24
<< metal1 >>
rect -40 28 -37 37
rect -36 25 -12 28
rect -8 25 16 28
rect 20 25 43 28
rect 47 25 71 28
rect -19 18 5 21
rect 9 18 33 21
rect 37 18 60 21
rect 64 18 88 21
rect -48 8 -35 11
rect -48 -1 -6 2
rect -48 -9 22 -6
rect -48 -19 48 -16
rect -48 -27 76 -24
rect 89 -33 92 18
rect -40 -46 -37 -43
<< labels >>
rlabel metal1 -39 34 -39 34 5 vdd!
rlabel metal1 -39 -44 -39 -44 1 gnd!
rlabel metal1 91 -11 91 -11 1 out
rlabel metal1 -47 10 -47 10 3 in1
rlabel metal1 -46 0 -46 0 3 in2
rlabel metal1 -47 -8 -47 -8 3 in3
rlabel metal1 -47 -18 -47 -18 3 in4
rlabel metal1 -46 -26 -46 -26 3 in5
<< end >>
