magic
tech scmos
timestamp 1699292645
<< nwell >>
rect -74 5 82 47
rect 96 7 134 46
<< ntransistor >>
rect -48 -31 -46 -5
rect -9 -31 -7 -5
rect 30 -31 32 -5
rect 63 -31 65 -5
rect 114 -29 116 -7
<< ptransistor >>
rect -48 13 -46 39
rect -9 13 -7 39
rect 30 13 32 39
rect 63 13 65 39
rect 114 15 116 37
<< ndiffusion >>
rect -60 -22 -48 -5
rect -56 -26 -48 -22
rect -60 -31 -48 -26
rect -46 -22 -29 -5
rect -46 -26 -38 -22
rect -34 -26 -29 -22
rect -46 -31 -29 -26
rect -23 -21 -9 -5
rect -23 -25 -21 -21
rect -17 -25 -9 -21
rect -23 -31 -9 -25
rect -7 -20 8 -5
rect -7 -24 3 -20
rect 7 -24 8 -20
rect -7 -31 8 -24
rect 12 -20 30 -5
rect 12 -24 17 -20
rect 21 -24 30 -20
rect 12 -31 30 -24
rect 32 -19 43 -5
rect 32 -23 37 -19
rect 41 -23 43 -19
rect 32 -31 43 -23
rect 48 -18 63 -5
rect 48 -22 50 -18
rect 54 -22 63 -18
rect 48 -31 63 -22
rect 65 -17 79 -5
rect 65 -21 70 -17
rect 74 -21 79 -17
rect 65 -31 79 -21
rect 106 -13 114 -7
rect 110 -17 114 -13
rect 106 -29 114 -17
rect 116 -14 129 -7
rect 116 -18 125 -14
rect 116 -29 129 -18
<< pdiffusion >>
rect -61 33 -48 39
rect -61 29 -58 33
rect -54 29 -48 33
rect -61 13 -48 29
rect -46 13 -9 39
rect -7 13 30 39
rect 32 13 63 39
rect 65 35 68 39
rect 65 13 72 35
rect 104 35 114 37
rect 108 31 114 35
rect 104 15 114 31
rect 116 29 127 37
rect 116 25 123 29
rect 116 15 127 25
<< ndcontact >>
rect -60 -26 -56 -22
rect -38 -26 -34 -22
rect -21 -25 -17 -21
rect 3 -24 7 -20
rect 17 -24 21 -20
rect 37 -23 41 -19
rect 50 -22 54 -18
rect 70 -21 74 -17
rect 106 -17 110 -13
rect 125 -18 129 -14
<< pdcontact >>
rect -58 29 -54 33
rect 68 35 72 39
rect 104 31 108 35
rect 123 25 127 29
<< polysilicon >>
rect -48 39 -46 42
rect -9 39 -7 42
rect 30 39 32 42
rect 63 39 65 42
rect 114 37 116 40
rect -48 -5 -46 13
rect -9 -5 -7 13
rect 30 -5 32 13
rect 63 -5 65 13
rect 114 -7 116 15
rect -48 -34 -46 -31
rect -9 -34 -7 -31
rect 30 -34 32 -31
rect 63 -34 65 -31
rect 114 -32 116 -29
<< polycontact >>
rect 110 0 114 4
<< metal1 >>
rect 72 35 89 38
rect 86 34 89 35
rect 86 31 104 34
rect -59 4 -55 29
rect -59 0 110 4
rect -59 -22 -55 0
rect 86 -17 106 -14
rect 124 -14 128 25
rect 74 -20 89 -17
rect -59 -38 -56 -26
rect -21 -37 -18 -25
rect 18 -34 21 -24
rect 51 -34 54 -22
rect 18 -37 54 -34
rect -21 -38 21 -37
rect -59 -41 21 -38
<< labels >>
rlabel metal1 126 2 126 2 1 out
rlabel metal1 89 32 89 32 1 vdd!
rlabel metal1 86 -19 86 -19 1 gnd!
rlabel ndcontact -36 -24 -36 -24 1 gnd!
rlabel ndcontact 5 -22 5 -22 1 gnd!
rlabel ndcontact 40 -21 40 -21 1 gnd!
rlabel polysilicon -47 40 -47 40 1 in1
rlabel polysilicon -8 41 -8 41 1 in2
rlabel polysilicon 31 41 31 41 1 in3
rlabel polysilicon 64 40 64 40 1 in4
<< end >>
