magic
tech scmos
timestamp 1700592115
<< nwell >>
rect -158 4 -126 22
rect -120 4 -87 22
rect -69 5 -6 28
rect -68 -16 -6 5
rect 18 4 50 22
rect 56 4 89 22
rect 107 5 170 28
rect 108 -16 170 5
rect 200 4 232 22
rect 238 4 271 22
rect 289 5 352 28
rect 290 -16 352 5
rect 382 4 414 22
rect 420 4 453 22
rect 471 5 534 28
rect 472 -16 534 5
rect -166 -102 -6 -80
rect 28 -101 164 -79
rect 202 -80 293 -76
rect 202 -98 314 -80
rect 293 -100 314 -98
rect 395 -104 459 -84
rect -120 -158 17 -136
<< ntransistor >>
rect -144 -12 -142 -6
rect -104 -12 -102 -6
rect 32 -12 34 -6
rect 72 -12 74 -6
rect 214 -12 216 -6
rect 254 -12 256 -6
rect 396 -12 398 -6
rect 436 -12 438 -6
rect -52 -30 -50 -23
rect -27 -30 -25 -23
rect 124 -30 126 -23
rect 149 -30 151 -23
rect 306 -30 308 -23
rect 331 -30 333 -23
rect 488 -30 490 -23
rect 513 -30 515 -23
rect -52 -47 -50 -39
rect -27 -47 -25 -39
rect 124 -47 126 -39
rect 149 -47 151 -39
rect 306 -47 308 -39
rect 331 -47 333 -39
rect 488 -47 490 -39
rect 513 -47 515 -39
rect -153 -123 -151 -113
rect -127 -123 -125 -113
rect -96 -123 -94 -113
rect -70 -123 -68 -113
rect -43 -123 -41 -113
rect -20 -119 -18 -114
rect 43 -122 45 -112
rect 74 -122 76 -112
rect 100 -122 102 -112
rect 127 -122 129 -112
rect 150 -118 152 -113
rect 217 -119 219 -109
rect 248 -119 250 -109
rect 274 -119 276 -109
rect 301 -114 303 -106
rect 406 -118 408 -110
rect 416 -118 418 -110
rect 443 -118 445 -110
rect -103 -179 -101 -169
rect -72 -179 -70 -169
rect -46 -179 -44 -169
rect -19 -179 -17 -169
rect 4 -175 6 -170
<< ptransistor >>
rect -144 10 -142 16
rect -104 10 -102 16
rect -52 15 -50 21
rect -28 15 -26 21
rect 32 10 34 16
rect 72 10 74 16
rect 124 15 126 21
rect 148 15 150 21
rect -51 -7 -49 0
rect -27 -7 -25 0
rect 214 10 216 16
rect 254 10 256 16
rect 306 15 308 21
rect 330 15 334 21
rect 125 -6 127 0
rect 149 -6 151 0
rect 396 10 398 16
rect 436 10 438 16
rect 488 15 490 21
rect 512 15 516 21
rect 307 -6 309 0
rect 330 -6 332 0
rect 489 -6 491 0
rect 512 -6 514 0
rect -153 -96 -151 -86
rect -127 -96 -125 -86
rect -96 -96 -94 -86
rect -70 -96 -68 -86
rect -43 -96 -41 -88
rect -20 -96 -18 -92
rect 43 -95 45 -85
rect 74 -95 76 -85
rect 100 -95 102 -85
rect 127 -95 129 -87
rect 150 -95 152 -91
rect 217 -92 219 -82
rect 248 -92 250 -82
rect 274 -92 276 -82
rect 301 -92 303 -86
rect 406 -98 408 -90
rect 416 -98 418 -90
rect 443 -98 445 -90
rect -103 -152 -101 -142
rect -72 -152 -70 -142
rect -46 -152 -44 -142
rect -19 -152 -17 -144
rect 4 -152 6 -148
<< ndiffusion >>
rect -148 -10 -144 -6
rect -152 -12 -144 -10
rect -142 -10 -137 -6
rect -142 -12 -133 -10
rect -109 -10 -104 -6
rect -113 -12 -104 -10
rect -102 -10 -98 -6
rect -102 -12 -94 -10
rect 29 -11 32 -6
rect 24 -12 32 -11
rect 34 -10 39 -6
rect 34 -12 43 -10
rect 67 -10 72 -6
rect 63 -12 72 -10
rect 74 -10 78 -6
rect 74 -12 82 -10
rect 211 -11 214 -6
rect 206 -12 214 -11
rect 216 -10 221 -6
rect 216 -12 225 -10
rect 249 -10 254 -6
rect 245 -12 254 -10
rect 256 -10 260 -6
rect 256 -12 264 -10
rect 393 -11 396 -6
rect 388 -12 396 -11
rect 398 -10 403 -6
rect 398 -12 407 -10
rect 431 -10 436 -6
rect 427 -12 436 -10
rect 438 -10 442 -6
rect 438 -12 446 -10
rect -42 -23 -37 -22
rect -61 -26 -52 -23
rect -57 -30 -52 -26
rect -50 -30 -27 -23
rect -25 -26 -11 -23
rect -25 -30 -15 -26
rect 115 -26 124 -23
rect 119 -30 124 -26
rect 126 -27 134 -23
rect 139 -27 149 -23
rect 126 -30 149 -27
rect 151 -26 165 -23
rect 151 -30 161 -26
rect 297 -26 306 -23
rect 301 -30 306 -26
rect 308 -27 316 -23
rect 321 -27 331 -23
rect 308 -30 331 -27
rect 333 -26 347 -23
rect 333 -30 343 -26
rect 479 -26 488 -23
rect 483 -30 488 -26
rect 490 -27 498 -23
rect 503 -27 513 -23
rect 490 -30 513 -27
rect 515 -26 529 -23
rect 515 -30 525 -26
rect -57 -43 -52 -39
rect -61 -47 -52 -43
rect -50 -43 -41 -39
rect -37 -43 -27 -39
rect -50 -47 -27 -43
rect -25 -43 -15 -39
rect -25 -47 -11 -43
rect 119 -43 124 -39
rect 115 -47 124 -43
rect 126 -43 135 -39
rect 139 -43 149 -39
rect 126 -47 149 -43
rect 151 -43 161 -39
rect 151 -47 165 -43
rect 301 -43 306 -39
rect 297 -47 306 -43
rect 308 -43 317 -39
rect 321 -43 331 -39
rect 308 -47 331 -43
rect 333 -43 343 -39
rect 333 -47 347 -43
rect 483 -43 488 -39
rect 479 -47 488 -43
rect 490 -43 499 -39
rect 503 -43 513 -39
rect 490 -47 513 -43
rect 515 -43 525 -39
rect 515 -47 529 -43
rect -161 -119 -153 -113
rect -157 -123 -153 -119
rect -151 -123 -127 -113
rect -125 -123 -96 -113
rect -94 -123 -70 -113
rect -68 -123 -43 -113
rect -41 -117 -38 -113
rect -41 -123 -34 -117
rect -22 -118 -20 -114
rect -24 -119 -20 -118
rect -18 -118 -16 -114
rect 38 -116 43 -112
rect -18 -119 -13 -118
rect 34 -122 43 -116
rect 45 -122 74 -112
rect 76 -122 100 -112
rect 102 -122 127 -112
rect 129 -116 132 -112
rect 212 -113 217 -109
rect 129 -122 136 -116
rect 148 -117 150 -113
rect 146 -118 150 -117
rect 152 -117 154 -113
rect 152 -118 157 -117
rect 208 -119 217 -113
rect 219 -119 248 -109
rect 250 -119 274 -109
rect 276 -113 282 -109
rect 276 -119 286 -113
rect 300 -110 301 -106
rect 296 -114 301 -110
rect 303 -110 305 -106
rect 303 -114 309 -110
rect 405 -114 406 -110
rect 401 -118 406 -114
rect 408 -118 416 -110
rect 418 -114 421 -110
rect 418 -118 425 -114
rect 442 -114 443 -110
rect 438 -118 443 -114
rect 445 -114 447 -110
rect 445 -118 451 -114
rect -108 -173 -103 -169
rect -112 -179 -103 -173
rect -101 -179 -72 -169
rect -70 -179 -46 -169
rect -44 -179 -19 -169
rect -17 -173 -14 -169
rect -17 -179 -10 -173
rect 2 -174 4 -170
rect 0 -175 4 -174
rect 6 -174 8 -170
rect 6 -175 11 -174
<< pdiffusion >>
rect -59 17 -52 21
rect -151 15 -144 16
rect -146 10 -144 15
rect -142 14 -132 16
rect -142 10 -136 14
rect -114 14 -104 16
rect -110 10 -104 14
rect -102 14 -95 16
rect -63 15 -52 17
rect -50 19 -28 21
rect -50 15 -42 19
rect -38 15 -28 19
rect -26 17 -17 21
rect -26 15 -13 17
rect 117 17 124 21
rect 25 15 32 16
rect -102 10 -99 14
rect 30 10 32 15
rect 34 14 44 16
rect 34 10 40 14
rect 62 14 72 16
rect 66 10 72 14
rect 74 14 81 16
rect 113 15 124 17
rect 126 19 148 21
rect 126 15 134 19
rect 138 15 148 19
rect 150 17 159 21
rect 150 15 163 17
rect 299 17 306 21
rect 207 15 214 16
rect 74 10 77 14
rect -58 -4 -51 0
rect -62 -7 -51 -4
rect -49 -3 -27 0
rect -49 -7 -41 -3
rect -37 -7 -27 -3
rect -25 -4 -16 0
rect -25 -7 -12 -4
rect 212 10 214 15
rect 216 14 226 16
rect 216 10 222 14
rect 244 14 254 16
rect 248 10 254 14
rect 256 14 263 16
rect 295 15 306 17
rect 308 19 330 21
rect 308 15 316 19
rect 320 15 330 19
rect 334 17 341 21
rect 334 15 345 17
rect 481 17 488 21
rect 389 15 396 16
rect 256 10 259 14
rect 118 -4 125 0
rect 114 -6 125 -4
rect 127 -2 149 0
rect 127 -6 135 -2
rect 139 -6 149 -2
rect 151 -4 160 0
rect 151 -6 164 -4
rect 394 10 396 15
rect 398 14 408 16
rect 398 10 404 14
rect 426 14 436 16
rect 430 10 436 14
rect 438 14 445 16
rect 477 15 488 17
rect 490 19 512 21
rect 490 15 498 19
rect 502 15 512 19
rect 516 17 523 21
rect 516 15 527 17
rect 438 10 441 14
rect 300 -4 307 0
rect 296 -6 307 -4
rect 309 -2 330 0
rect 309 -6 317 -2
rect 321 -6 330 -2
rect 332 -4 342 0
rect 332 -6 346 -4
rect 482 -4 489 0
rect 478 -6 489 -4
rect 491 -2 512 0
rect 491 -6 499 -2
rect 503 -6 512 -2
rect 514 -4 524 0
rect 514 -6 528 -4
rect -159 -92 -153 -86
rect -155 -96 -153 -92
rect -151 -92 -144 -86
rect -151 -96 -148 -92
rect -136 -92 -127 -86
rect -132 -96 -127 -92
rect -125 -92 -117 -86
rect -125 -96 -121 -92
rect -106 -92 -96 -86
rect -102 -96 -96 -92
rect -94 -92 -84 -86
rect -94 -96 -88 -92
rect -79 -92 -70 -86
rect -75 -96 -70 -92
rect -68 -92 -58 -86
rect -68 -96 -62 -92
rect -50 -92 -43 -88
rect -46 -96 -43 -92
rect -41 -92 -32 -88
rect 34 -91 43 -85
rect -41 -96 -36 -92
rect -22 -96 -20 -92
rect -18 -96 -17 -92
rect 38 -95 43 -91
rect 45 -91 53 -85
rect 45 -95 49 -91
rect 64 -91 74 -85
rect 68 -95 74 -91
rect 76 -91 86 -85
rect 76 -95 82 -91
rect 91 -91 100 -85
rect 95 -95 100 -91
rect 102 -91 112 -85
rect 102 -95 108 -91
rect 120 -91 127 -87
rect 124 -95 127 -91
rect 129 -91 138 -87
rect 208 -88 217 -82
rect 129 -95 134 -91
rect 148 -95 150 -91
rect 152 -95 153 -91
rect 212 -92 217 -88
rect 219 -88 227 -82
rect 219 -92 223 -88
rect 238 -88 248 -82
rect 242 -92 248 -88
rect 250 -88 260 -82
rect 250 -92 256 -88
rect 265 -88 274 -82
rect 269 -92 274 -88
rect 276 -88 286 -82
rect 276 -92 282 -88
rect 300 -90 301 -86
rect 296 -92 301 -90
rect 303 -88 308 -86
rect 303 -92 304 -88
rect 401 -94 406 -90
rect 405 -98 406 -94
rect 408 -94 416 -90
rect 408 -98 410 -94
rect 414 -98 416 -94
rect 418 -94 425 -90
rect 418 -98 421 -94
rect 438 -94 443 -90
rect 442 -98 443 -94
rect 445 -94 450 -90
rect 445 -98 446 -94
rect -112 -148 -103 -142
rect -108 -152 -103 -148
rect -101 -148 -93 -142
rect -101 -152 -97 -148
rect -82 -148 -72 -142
rect -78 -152 -72 -148
rect -70 -148 -60 -142
rect -70 -152 -64 -148
rect -55 -148 -46 -142
rect -51 -152 -46 -148
rect -44 -148 -34 -142
rect -44 -152 -38 -148
rect -26 -148 -19 -144
rect -22 -152 -19 -148
rect -17 -148 -8 -144
rect -17 -152 -12 -148
rect 2 -152 4 -148
rect 6 -152 7 -148
<< ndcontact >>
rect -152 -10 -148 -6
rect -137 -10 -133 -6
rect -113 -10 -109 -6
rect -98 -10 -94 -6
rect 39 -10 43 -6
rect 63 -10 67 -6
rect 78 -10 82 -6
rect 221 -10 225 -6
rect 245 -10 249 -6
rect 260 -10 264 -6
rect 403 -10 407 -6
rect 427 -10 431 -6
rect 442 -10 446 -6
rect -61 -30 -57 -26
rect -15 -30 -11 -26
rect 115 -30 119 -26
rect 134 -27 139 -22
rect 161 -30 165 -26
rect 297 -30 301 -26
rect 316 -27 321 -22
rect 343 -30 347 -26
rect 479 -30 483 -26
rect 498 -27 503 -22
rect 525 -30 529 -26
rect -61 -43 -57 -39
rect -41 -43 -37 -39
rect -15 -43 -11 -39
rect 115 -43 119 -39
rect 135 -43 139 -39
rect 161 -43 165 -39
rect 297 -43 301 -39
rect 317 -43 321 -39
rect 343 -43 347 -39
rect 479 -43 483 -39
rect 499 -43 503 -39
rect 525 -43 529 -39
rect -161 -123 -157 -119
rect -38 -117 -34 -113
rect -26 -118 -22 -114
rect -16 -118 -12 -114
rect 34 -116 38 -112
rect 132 -116 136 -112
rect 208 -113 212 -109
rect 144 -117 148 -113
rect 154 -117 158 -113
rect 282 -113 286 -109
rect 296 -110 300 -106
rect 305 -110 309 -106
rect 401 -114 405 -110
rect 421 -114 425 -110
rect 438 -114 442 -110
rect 447 -114 451 -110
rect -112 -173 -108 -169
rect -14 -173 -10 -169
rect -2 -174 2 -170
rect 8 -174 12 -170
<< pdcontact >>
rect -63 17 -59 21
rect -136 10 -132 14
rect -114 10 -110 14
rect -42 15 -38 19
rect -17 17 -13 21
rect 113 17 117 21
rect -99 10 -95 14
rect 40 10 44 14
rect 62 10 66 14
rect 134 15 138 19
rect 159 17 163 21
rect 295 17 299 21
rect 77 10 81 14
rect -62 -4 -58 0
rect -41 -7 -37 -3
rect -16 -4 -12 0
rect 222 10 226 14
rect 244 10 248 14
rect 316 15 320 19
rect 341 17 345 21
rect 477 17 481 21
rect 259 10 263 14
rect 114 -4 118 0
rect 135 -6 139 -2
rect 160 -4 164 0
rect 404 10 408 14
rect 426 10 430 14
rect 498 15 502 19
rect 523 17 527 21
rect 441 10 445 14
rect 296 -4 300 0
rect 317 -6 321 -2
rect 342 -4 346 0
rect 478 -4 482 0
rect 499 -6 503 -2
rect 524 -4 528 0
rect -159 -96 -155 -92
rect -148 -96 -144 -92
rect -136 -96 -132 -92
rect -121 -96 -117 -92
rect -106 -96 -102 -92
rect -88 -96 -84 -92
rect -79 -96 -75 -92
rect -62 -96 -58 -92
rect -50 -96 -46 -92
rect -36 -96 -32 -92
rect -26 -96 -22 -92
rect -17 -96 -13 -92
rect 34 -95 38 -91
rect 49 -95 53 -91
rect 64 -95 68 -91
rect 82 -95 86 -91
rect 91 -95 95 -91
rect 108 -95 112 -91
rect 120 -95 124 -91
rect 134 -95 138 -91
rect 144 -95 148 -91
rect 153 -95 157 -91
rect 208 -92 212 -88
rect 223 -92 227 -88
rect 238 -92 242 -88
rect 256 -92 260 -88
rect 265 -92 269 -88
rect 282 -92 286 -88
rect 296 -90 300 -86
rect 304 -92 308 -88
rect 401 -98 405 -94
rect 410 -98 414 -94
rect 421 -98 425 -94
rect 438 -98 442 -94
rect 446 -98 450 -94
rect -112 -152 -108 -148
rect -97 -152 -93 -148
rect -82 -152 -78 -148
rect -64 -152 -60 -148
rect -55 -152 -51 -148
rect -38 -152 -34 -148
rect -26 -152 -22 -148
rect -12 -152 -8 -148
rect -2 -152 2 -148
rect 7 -152 11 -148
<< polysilicon >>
rect -52 21 -50 24
rect -28 21 -26 24
rect 124 21 126 24
rect 148 21 150 24
rect 306 21 308 24
rect 330 21 334 24
rect 488 21 490 24
rect 512 21 516 24
rect -144 16 -142 19
rect -104 16 -102 19
rect 32 16 34 19
rect 72 16 74 19
rect -52 14 -50 15
rect -28 14 -26 15
rect -144 -6 -142 10
rect -104 4 -102 10
rect -51 10 -50 14
rect -27 10 -26 14
rect 214 16 216 19
rect 254 16 256 19
rect 124 14 126 15
rect 148 14 150 15
rect -108 -1 -102 4
rect -51 0 -49 3
rect -27 0 -25 3
rect -104 -6 -102 -1
rect 32 -6 34 10
rect 72 3 74 10
rect 125 10 126 14
rect 149 10 150 14
rect 396 16 398 19
rect 436 16 438 19
rect 306 14 308 15
rect 67 -2 74 3
rect 125 0 127 3
rect 149 0 151 3
rect 72 -6 74 -2
rect 214 -6 216 10
rect 254 3 256 10
rect 307 10 308 14
rect 330 10 334 15
rect 488 14 490 15
rect 249 -2 256 3
rect 307 0 309 3
rect 330 0 332 3
rect 254 -6 256 -2
rect 396 -6 398 10
rect 436 3 438 10
rect 489 10 490 14
rect 512 10 516 15
rect 431 -2 438 3
rect 489 0 491 3
rect 512 0 514 3
rect 436 -6 438 -2
rect -144 -15 -142 -12
rect -104 -15 -102 -12
rect -51 -13 -49 -7
rect -27 -13 -25 -7
rect 32 -15 34 -12
rect 72 -15 74 -12
rect 125 -13 127 -6
rect 149 -13 151 -6
rect 214 -15 216 -12
rect 254 -15 256 -12
rect 307 -13 309 -6
rect 330 -13 332 -6
rect 396 -15 398 -12
rect 436 -15 438 -12
rect 489 -13 491 -6
rect 512 -13 514 -6
rect -52 -23 -50 -17
rect -27 -23 -25 -17
rect 124 -23 126 -17
rect 149 -23 151 -17
rect 306 -23 308 -17
rect 331 -23 333 -17
rect 488 -23 490 -17
rect 513 -23 515 -17
rect -52 -33 -50 -30
rect -27 -33 -25 -30
rect 124 -33 126 -30
rect 149 -33 151 -30
rect 306 -33 308 -30
rect 331 -33 333 -30
rect 488 -33 490 -30
rect 513 -33 515 -30
rect -52 -39 -50 -36
rect -27 -39 -25 -36
rect 124 -39 126 -36
rect 149 -39 151 -36
rect 306 -39 308 -36
rect 331 -39 333 -36
rect 488 -39 490 -36
rect 513 -39 515 -36
rect -52 -57 -50 -47
rect -27 -54 -25 -47
rect 124 -56 126 -47
rect 149 -54 151 -47
rect 306 -54 308 -47
rect 331 -54 333 -47
rect 488 -54 490 -47
rect 513 -54 515 -47
rect -153 -86 -151 -79
rect -127 -86 -125 -79
rect -96 -86 -94 -79
rect -70 -86 -68 -79
rect -43 -88 -41 -79
rect 43 -85 45 -70
rect 100 -70 102 -68
rect 74 -85 76 -71
rect 100 -85 102 -75
rect -20 -92 -18 -89
rect 127 -87 129 -73
rect 217 -82 219 -69
rect 248 -82 250 -65
rect 274 -82 276 -73
rect 407 -79 408 -76
rect 150 -91 152 -88
rect 301 -86 303 -83
rect 406 -90 408 -79
rect 416 -90 418 -75
rect 443 -90 445 -87
rect -153 -113 -151 -96
rect -127 -113 -125 -96
rect -96 -113 -94 -96
rect -70 -113 -68 -96
rect -43 -113 -41 -96
rect -20 -114 -18 -96
rect 43 -112 45 -95
rect 74 -112 76 -95
rect 100 -112 102 -95
rect 127 -112 129 -95
rect -20 -122 -18 -119
rect 150 -113 152 -95
rect 217 -109 219 -92
rect 248 -109 250 -92
rect 274 -109 276 -92
rect 301 -106 303 -92
rect 150 -121 152 -118
rect 406 -110 408 -98
rect 416 -110 418 -98
rect 443 -110 445 -98
rect 301 -118 303 -114
rect 217 -122 219 -119
rect 248 -122 250 -119
rect 274 -122 276 -119
rect 406 -121 408 -118
rect 416 -121 418 -118
rect 443 -121 445 -118
rect -153 -127 -151 -123
rect -127 -126 -125 -123
rect -96 -126 -94 -123
rect -70 -126 -68 -123
rect -43 -126 -41 -123
rect 43 -125 45 -122
rect 74 -125 76 -122
rect 100 -125 102 -122
rect 127 -125 129 -122
rect -71 -138 -70 -134
rect -103 -142 -101 -138
rect -72 -142 -70 -138
rect -46 -142 -44 -138
rect -19 -144 -17 -139
rect 4 -148 6 -145
rect -103 -169 -101 -152
rect -72 -169 -70 -152
rect -46 -169 -44 -152
rect -19 -169 -17 -152
rect 4 -170 6 -152
rect 4 -178 6 -175
rect -103 -182 -101 -179
rect -72 -182 -70 -179
rect -46 -182 -44 -179
rect -19 -182 -17 -179
<< polycontact >>
rect 332 -12 336 -8
rect 514 -12 518 -8
rect 42 -70 47 -65
rect -151 -82 -146 -77
rect -125 -82 -120 -77
rect -94 -82 -89 -77
rect -68 -82 -63 -77
rect -41 -83 -36 -78
rect 74 -71 79 -66
rect 216 -69 221 -64
rect 100 -75 105 -70
rect 129 -77 134 -72
rect 250 -69 255 -64
rect 276 -76 281 -71
rect 402 -79 407 -74
rect 418 -78 423 -73
rect -24 -106 -20 -102
rect 146 -105 150 -101
rect 297 -103 301 -99
rect 439 -106 443 -102
rect -106 -138 -101 -133
rect -76 -138 -71 -133
rect -49 -138 -44 -133
rect 0 -162 4 -158
<< metal1 >>
rect -63 25 55 28
rect -63 23 -60 25
rect -124 22 -60 23
rect -172 21 -60 22
rect -17 21 -14 25
rect 51 23 55 25
rect 113 25 238 28
rect 113 23 116 25
rect 51 21 116 23
rect 159 21 162 25
rect 170 24 238 25
rect 234 23 238 24
rect 295 25 419 28
rect 295 23 298 25
rect 234 21 298 23
rect 341 21 344 25
rect 416 23 419 25
rect 477 25 534 28
rect 477 23 480 25
rect 416 21 480 23
rect 523 21 526 25
rect -172 20 -63 21
rect -172 19 -121 20
rect -172 -93 -169 19
rect -124 13 -121 19
rect 52 20 113 21
rect -132 10 -114 13
rect -151 -6 -148 10
rect -98 0 -95 10
rect -42 6 -39 15
rect 52 13 55 20
rect 234 20 295 21
rect 44 10 62 13
rect -62 3 -13 6
rect -62 0 -59 3
rect -16 0 -13 3
rect -98 -3 -83 0
rect -98 -6 -95 -3
rect -133 -10 -113 -7
rect -86 -9 -83 -3
rect 25 -6 28 10
rect 78 0 81 10
rect 134 6 137 15
rect 234 13 237 20
rect 416 20 477 21
rect 226 10 244 13
rect 114 3 163 6
rect 114 0 117 3
rect 160 0 163 3
rect 78 -3 93 0
rect 78 -6 81 -3
rect -125 -19 -122 -10
rect -86 -12 -56 -9
rect -125 -22 -74 -19
rect -41 -22 -38 -7
rect 43 -10 63 -7
rect 90 -9 93 -3
rect 207 -6 210 10
rect 260 0 263 10
rect 316 6 319 15
rect 416 13 419 20
rect 408 10 426 13
rect 296 3 345 6
rect 296 0 299 3
rect 342 0 345 3
rect 260 -3 275 0
rect 260 -6 263 -3
rect 51 -19 54 -10
rect 90 -12 120 -9
rect 51 -22 102 -19
rect 135 -22 138 -6
rect 225 -10 245 -7
rect 272 -9 275 -3
rect 389 -6 392 10
rect 442 0 445 10
rect 498 6 501 15
rect 478 3 527 6
rect 478 0 481 3
rect 524 0 527 3
rect 442 -3 457 0
rect 442 -6 445 -3
rect 233 -19 236 -10
rect 272 -12 302 -9
rect 233 -22 284 -19
rect 317 -22 320 -6
rect 349 -7 352 -6
rect 336 -11 347 -8
rect 407 -10 427 -7
rect 454 -9 457 -3
rect 389 -12 392 -11
rect 415 -19 418 -10
rect 454 -12 484 -9
rect 415 -22 466 -19
rect 499 -22 502 -6
rect 531 -7 534 -6
rect 518 -11 529 -8
rect -77 -47 -74 -22
rect -61 -39 -58 -30
rect -14 -39 -11 -30
rect -63 -47 -46 -46
rect -41 -47 -38 -43
rect -77 -49 -38 -47
rect -77 -50 -60 -49
rect -49 -50 -38 -49
rect 99 -47 102 -22
rect 115 -39 118 -30
rect 162 -39 165 -30
rect 113 -47 130 -46
rect 135 -47 138 -43
rect 99 -49 138 -47
rect 281 -47 284 -22
rect 297 -39 300 -30
rect 344 -39 347 -30
rect 295 -47 312 -46
rect 317 -47 320 -43
rect 281 -49 320 -47
rect 463 -47 466 -22
rect 479 -39 482 -30
rect 526 -39 529 -30
rect 499 -47 502 -43
rect 99 -50 116 -49
rect 127 -50 138 -49
rect -41 -58 -38 -50
rect 135 -57 138 -50
rect 281 -50 298 -49
rect 309 -50 320 -49
rect 317 -57 320 -50
rect 463 -50 502 -47
rect 362 -57 365 -56
rect 135 -58 253 -57
rect 317 -58 435 -57
rect -41 -60 74 -58
rect 132 -59 264 -58
rect 315 -59 441 -58
rect 132 -60 292 -59
rect 309 -60 441 -59
rect -41 -61 292 -60
rect 299 -61 441 -60
rect 71 -63 135 -61
rect 261 -62 318 -61
rect 289 -63 312 -62
rect 289 -64 309 -63
rect 438 -67 441 -61
rect 499 -67 502 -50
rect 438 -70 502 -67
rect -68 -77 -64 -75
rect 281 -76 288 -73
rect 402 -74 406 -72
rect 423 -78 426 -75
rect 362 -82 365 -81
rect 208 -85 426 -82
rect 34 -86 211 -85
rect -159 -88 211 -86
rect 238 -88 242 -85
rect 266 -88 269 -85
rect 296 -86 300 -85
rect -159 -89 37 -88
rect -159 -92 -156 -89
rect -136 -92 -133 -89
rect -106 -92 -102 -89
rect -78 -92 -75 -89
rect -50 -92 -47 -89
rect -26 -92 -23 -89
rect 34 -91 37 -89
rect 64 -91 68 -88
rect 92 -91 95 -88
rect 120 -91 123 -88
rect 144 -91 147 -88
rect -172 -96 -159 -93
rect -172 -143 -168 -96
rect -147 -103 -144 -96
rect -121 -103 -118 -96
rect -87 -103 -84 -96
rect -61 -103 -58 -96
rect -35 -103 -32 -96
rect -147 -106 -24 -103
rect -38 -113 -35 -106
rect -16 -114 -13 -96
rect 49 -102 52 -95
rect 83 -102 86 -95
rect 109 -102 112 -95
rect 135 -102 138 -95
rect 49 -105 146 -102
rect 132 -112 135 -105
rect 154 -113 157 -95
rect 223 -99 226 -92
rect 257 -99 260 -92
rect 283 -99 286 -92
rect 223 -102 297 -99
rect 283 -109 286 -102
rect 305 -106 308 -92
rect 401 -94 404 -85
rect 422 -94 426 -85
rect 425 -95 426 -94
rect 425 -98 438 -95
rect 411 -104 414 -98
rect 421 -104 439 -103
rect 411 -106 439 -104
rect 411 -107 424 -106
rect 421 -110 424 -107
rect 447 -110 450 -98
rect -161 -128 -158 -123
rect -112 -128 -95 -127
rect -82 -128 -65 -127
rect -55 -128 -38 -127
rect -26 -128 -23 -118
rect 34 -127 37 -116
rect 144 -127 147 -117
rect 208 -124 211 -113
rect 296 -124 299 -110
rect 401 -122 404 -114
rect 438 -121 441 -114
rect 499 -121 502 -70
rect 438 -122 502 -121
rect 398 -124 502 -122
rect 206 -125 502 -124
rect 206 -127 404 -125
rect 31 -128 209 -127
rect -161 -130 209 -128
rect -161 -131 -109 -130
rect -98 -131 -79 -130
rect -68 -131 -52 -130
rect -41 -131 34 -130
rect -71 -137 -70 -134
rect -112 -143 12 -142
rect -172 -145 12 -143
rect -172 -146 -109 -145
rect -112 -148 -109 -146
rect -82 -148 -78 -145
rect -54 -148 -51 -145
rect -26 -148 -23 -145
rect -2 -148 1 -145
rect -97 -159 -94 -152
rect -63 -159 -60 -152
rect -37 -159 -34 -152
rect -11 -159 -8 -152
rect -97 -162 0 -159
rect -14 -169 -11 -162
rect 8 -170 11 -152
rect -112 -185 -109 -173
rect -2 -184 1 -174
rect 21 -184 25 -131
rect -2 -185 25 -184
rect -112 -188 25 -185
<< m2contact >>
rect 347 -12 352 -7
rect 529 -12 534 -7
<< pm12contact >>
rect -142 -2 -137 3
rect -56 9 -51 14
rect -32 9 -27 14
rect 34 -2 39 3
rect 120 9 125 14
rect 144 9 149 14
rect -56 -13 -51 -8
rect -57 -22 -52 -17
rect -25 -13 -20 -8
rect 216 -2 221 3
rect 302 9 307 14
rect 325 9 330 14
rect -25 -22 -20 -17
rect 120 -13 125 -8
rect 119 -22 124 -17
rect 151 -12 156 -7
rect 398 -2 403 3
rect 484 9 489 14
rect 507 9 512 14
rect 151 -22 156 -17
rect 302 -13 307 -8
rect 301 -22 306 -17
rect 333 -22 338 -17
rect 484 -13 489 -8
rect 483 -22 488 -17
rect 515 -22 520 -17
rect -57 -57 -52 -52
rect -25 -55 -20 -50
rect 119 -57 124 -52
rect 151 -54 156 -49
rect 301 -57 306 -52
rect 333 -54 338 -49
rect 484 -59 490 -54
rect 515 -54 520 -49
rect -19 -139 -14 -134
<< pdm12contact >>
rect -151 10 -146 15
rect 25 10 30 15
rect 207 10 212 15
rect 389 10 394 15
<< ndm12contact >>
rect 24 -11 29 -6
rect 206 -11 211 -6
rect 388 -11 393 -6
<< metal2 >>
rect -163 32 -6 35
rect -163 3 -160 32
rect -151 25 -29 28
rect -151 15 -148 25
rect -32 14 -29 25
rect -66 10 -56 13
rect -163 0 -142 3
rect -66 3 -63 10
rect -103 0 -63 3
rect -151 -23 -148 -10
rect -66 -18 -63 0
rect -51 -13 -29 -10
rect -9 -10 -6 32
rect 13 32 170 35
rect 13 3 16 32
rect 25 25 147 28
rect 25 15 28 25
rect 144 14 147 25
rect 110 10 120 13
rect 110 3 113 10
rect 13 0 34 3
rect 72 0 113 3
rect -20 -13 -6 -10
rect -32 -17 -29 -13
rect -66 -21 -57 -18
rect -32 -20 -25 -17
rect -146 -26 -79 -23
rect -82 -52 -79 -26
rect -82 -55 -57 -52
rect -9 -51 -6 -13
rect -20 -54 -6 -51
rect -2 -135 1 -20
rect 25 -23 28 -11
rect 110 -18 113 0
rect 125 -13 147 -10
rect 167 -9 170 32
rect 195 32 352 35
rect 195 3 198 32
rect 207 25 329 28
rect 207 15 210 25
rect 326 14 329 25
rect 292 10 302 13
rect 292 3 295 10
rect 195 0 216 3
rect 254 0 295 3
rect 156 -12 170 -9
rect 144 -17 147 -13
rect 110 -21 119 -18
rect 144 -20 151 -17
rect 25 -26 33 -23
rect 39 -26 97 -23
rect 94 -52 97 -26
rect 94 -55 119 -52
rect 167 -51 170 -12
rect 207 -23 210 -11
rect 292 -18 295 0
rect 349 -7 352 32
rect 377 32 534 35
rect 377 3 380 32
rect 389 25 511 28
rect 389 15 392 25
rect 508 14 511 25
rect 474 10 484 13
rect 474 3 477 10
rect 377 0 398 3
rect 436 0 477 3
rect 307 -13 329 -10
rect 326 -17 329 -13
rect 292 -21 301 -18
rect 326 -20 333 -17
rect 207 -26 215 -23
rect 221 -26 279 -23
rect 156 -54 170 -51
rect 276 -52 279 -26
rect 276 -55 301 -52
rect 349 -51 352 -12
rect 389 -23 392 -11
rect 474 -18 477 0
rect 531 -7 534 32
rect 489 -13 511 -10
rect 508 -17 511 -13
rect 474 -21 483 -18
rect 508 -20 515 -17
rect 389 -26 398 -23
rect 403 -26 461 -23
rect 338 -54 352 -51
rect 458 -54 461 -26
rect 531 -51 534 -12
rect 520 -54 534 -51
rect 458 -57 484 -54
rect -14 -138 1 -135
<< m3contact >>
rect -151 -28 -146 -23
rect -2 -20 3 -15
rect -151 -82 -146 -77
rect -125 -82 -120 -77
rect -94 -82 -89 -77
rect -68 -82 -63 -77
rect -41 -83 -36 -78
rect -106 -138 -101 -133
rect -76 -138 -71 -133
rect -49 -138 -44 -133
rect 33 -28 39 -22
rect 134 -27 139 -22
rect 215 -28 221 -22
rect 316 -27 321 -22
rect 398 -27 403 -22
rect 498 -27 503 -22
rect 42 -70 47 -65
rect 74 -71 79 -66
rect 216 -69 221 -64
rect 250 -69 255 -64
rect 100 -75 105 -70
rect 129 -77 134 -72
rect 276 -76 281 -71
rect 402 -79 407 -74
rect 418 -78 423 -73
<< m123contact >>
rect -108 -1 -103 4
rect 67 -2 72 3
rect -42 -27 -37 -22
rect 249 -2 254 3
rect 431 -2 436 3
<< metal3 >>
rect 355 40 358 41
rect 5 36 176 39
rect -125 -1 -108 2
rect -151 -77 -148 -28
rect -125 -77 -122 -1
rect 5 -8 9 36
rect 5 -11 13 -8
rect -41 -15 1 -14
rect -41 -17 -2 -15
rect -41 -22 -38 -17
rect 9 -24 13 -11
rect 5 -27 13 -24
rect 5 -63 9 -27
rect -94 -66 9 -63
rect 35 -66 38 -28
rect 68 -63 71 -2
rect 173 -14 176 36
rect 135 -17 176 -14
rect 191 37 358 40
rect 135 -22 138 -17
rect 191 -61 194 37
rect -94 -77 -91 -66
rect 35 -69 42 -66
rect 68 -66 79 -63
rect 102 -64 194 -61
rect 216 -64 219 -28
rect 250 -64 253 -2
rect 355 -14 358 37
rect 317 -17 358 -14
rect 372 36 540 39
rect 317 -22 320 -17
rect 102 -70 105 -64
rect -48 -74 -29 -71
rect -48 -75 -45 -74
rect -76 -77 -45 -75
rect -106 -81 -94 -78
rect -106 -133 -103 -81
rect -76 -78 -68 -77
rect -76 -133 -73 -78
rect -63 -78 -45 -77
rect -32 -75 -29 -74
rect -32 -78 105 -75
rect 134 -76 276 -73
rect 372 -73 375 36
rect 281 -76 375 -73
rect 399 -72 402 -27
rect 399 -74 406 -72
rect 399 -75 402 -74
rect -50 -83 -41 -82
rect 129 -82 132 -77
rect 432 -75 435 -2
rect 537 -14 540 36
rect 499 -17 540 -14
rect 499 -22 502 -17
rect 423 -78 435 -75
rect -36 -83 133 -82
rect -50 -85 133 -83
rect -50 -133 -47 -85
rect -71 -137 -70 -134
rect -50 -137 -49 -133
<< labels >>
rlabel polysilicon -103 0 -103 0 1 a0
rlabel polysilicon -144 0 -142 2 1 b0
rlabel pm12contact 36 1 36 1 1 b1
rlabel metal1 70 0 70 0 1 a1
rlabel pm12contact 219 1 219 1 1 b2
rlabel m123contact 251 1 251 1 1 a2
rlabel pm12contact 400 1 400 1 1 b3
rlabel m123contact 435 1 435 1 1 a3
rlabel metal3 -2 -15 -2 -15 1 w0
rlabel metal1 449 -105 449 -105 1 s3
rlabel metal1 305 -102 308 -100 1 s2
rlabel metal1 155 -103 155 -103 1 s1
rlabel metal1 -14 -105 -14 -105 1 s0
rlabel metal1 10 -160 10 -160 1 A_gr
rlabel metal1 -170 -46 -170 -46 3 vdd!
rlabel metal1 500 -82 500 -82 1 gnd!
rlabel m3contact 137 -24 137 -24 1 w1
rlabel m3contact 318 -24 318 -24 1 w2
rlabel metal3 500 -20 500 -20 1 w3
<< end >>
