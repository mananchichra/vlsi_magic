magic
tech scmos
timestamp 1701288896
<< nwell >>
rect 120 -314 123 -293
<< polysilicon >>
rect -370 35 -368 150
rect 243 112 247 114
rect 256 112 260 120
rect -442 -79 -440 -34
rect -409 -68 -407 -32
rect -370 -52 -368 -35
rect -409 -70 -384 -68
rect -442 -81 -401 -79
rect -403 -268 -401 -81
rect -386 -178 -384 -70
rect -331 -82 -329 -34
rect -386 -180 -362 -178
rect -403 -270 -275 -268
<< polycontact >>
rect -372 150 -367 154
rect 256 120 260 124
rect 243 114 247 118
rect -333 -86 -329 -82
rect -362 -181 -357 -177
rect -279 -274 -275 -270
<< metal1 >>
rect -209 283 -24 289
rect -216 277 -203 283
rect -216 267 -210 277
rect -280 261 -210 267
rect -30 266 -24 283
rect -280 245 -274 261
rect -30 260 17 266
rect -336 239 -274 245
rect -193 251 -180 254
rect -153 251 -122 254
rect -336 229 -330 239
rect -503 223 -330 229
rect -193 228 -190 251
rect -305 225 -233 228
rect -193 225 -145 228
rect -503 63 -497 223
rect -305 216 -302 225
rect -521 57 -497 63
rect -473 215 -302 216
rect -473 213 -321 215
rect -521 7 -515 57
rect -473 30 -470 213
rect -316 213 -302 215
rect -236 211 -233 225
rect -321 207 -316 210
rect -148 192 -145 225
rect -146 185 -143 186
rect -370 180 -338 183
rect -312 182 -284 185
rect -146 184 -142 185
rect -146 181 -128 184
rect -370 154 -366 180
rect -145 177 -143 178
rect -146 174 -135 177
rect -286 159 -282 162
rect -367 153 -366 154
rect -138 153 -135 174
rect -131 162 -128 181
rect -125 166 -122 251
rect 11 221 17 260
rect 11 215 145 221
rect 128 175 131 197
rect 139 190 145 215
rect 139 184 194 190
rect 70 171 96 174
rect 120 172 178 175
rect 70 169 74 171
rect 61 165 74 169
rect -131 159 -119 162
rect -138 150 -129 153
rect -132 87 -129 150
rect -132 84 140 87
rect -169 41 -158 44
rect -135 41 -126 44
rect -169 22 -166 41
rect -169 19 -144 22
rect -521 1 -504 7
rect -147 -5 -144 19
rect -129 9 -126 41
rect -129 6 -119 9
rect 66 5 80 8
rect 137 6 140 84
rect 77 2 104 5
rect 127 3 140 6
rect -125 1 -122 2
rect -154 -8 -144 -5
rect -134 -2 -122 1
rect -134 -12 -131 -2
rect -458 -13 -381 -12
rect -458 -15 -341 -13
rect -154 -15 -131 -12
rect -476 -72 -473 -15
rect -458 -21 -455 -15
rect -417 -21 -414 -15
rect -384 -16 -341 -15
rect -384 -21 -381 -16
rect -344 -23 -341 -16
rect -285 -21 -218 -17
rect -344 -26 -339 -23
rect -476 -75 -456 -72
rect -459 -115 -456 -75
rect -285 -83 -282 -21
rect -161 -23 -125 -20
rect -154 -30 -146 -27
rect -160 -44 -157 -42
rect -153 -68 -149 -30
rect -128 -64 -125 -23
rect 18 -23 21 -10
rect 108 -23 111 -9
rect 137 -20 140 3
rect 175 -14 178 172
rect 188 145 194 184
rect 188 139 262 145
rect 256 124 262 139
rect 260 123 262 124
rect 220 118 247 119
rect 220 114 243 118
rect 220 52 225 114
rect 228 99 238 103
rect 228 90 232 99
rect 266 85 278 89
rect 252 60 255 70
rect 252 57 337 60
rect 220 47 328 52
rect 200 2 203 6
rect 254 2 292 5
rect 293 -14 296 1
rect 175 -17 202 -14
rect 137 -23 195 -20
rect 18 -26 111 -23
rect 126 -32 193 -28
rect -329 -86 -319 -83
rect -292 -86 -282 -83
rect -194 -72 -149 -68
rect 126 -68 130 -32
rect 323 -35 328 47
rect 184 -37 199 -35
rect -194 -94 -190 -72
rect -128 -73 -125 -69
rect 13 -71 130 -68
rect 13 -73 16 -71
rect -128 -76 16 -73
rect -230 -98 -190 -94
rect 126 -83 130 -71
rect 165 -38 199 -37
rect 165 -40 187 -38
rect 262 -39 289 -36
rect 315 -40 329 -35
rect -459 -118 -429 -115
rect -432 -164 -429 -118
rect -230 -162 -226 -98
rect -168 -123 -159 -120
rect -136 -122 -127 -119
rect -168 -138 -165 -123
rect -168 -141 -149 -138
rect -432 -167 -407 -164
rect -410 -210 -407 -167
rect -231 -166 -226 -162
rect -152 -163 -149 -141
rect -130 -152 -127 -122
rect 126 -134 129 -83
rect 63 -138 95 -135
rect 119 -137 129 -134
rect 63 -152 67 -138
rect -130 -155 -119 -152
rect 63 -156 66 -152
rect -159 -166 -149 -163
rect -131 -162 -120 -159
rect -131 -169 -128 -162
rect -158 -172 -128 -169
rect -288 -174 -278 -173
rect -288 -177 -205 -174
rect -357 -180 -315 -177
rect -288 -179 -278 -177
rect -158 -178 -149 -175
rect -165 -192 -162 -188
rect -410 -213 -297 -210
rect -300 -342 -297 -213
rect -152 -230 -149 -178
rect 18 -183 21 -171
rect 100 -183 103 -147
rect 18 -186 103 -183
rect 165 -233 168 -40
rect 202 -66 205 -46
rect 292 -66 295 -48
rect 334 -66 337 57
rect 202 -69 337 -66
rect 202 -94 205 -69
rect 202 -97 219 -94
rect -147 -234 -52 -233
rect -40 -234 168 -233
rect -147 -235 168 -234
rect -152 -236 168 -235
rect -55 -237 -32 -236
rect -161 -272 -153 -269
rect -129 -271 -122 -268
rect -279 -298 -276 -274
rect -279 -301 -261 -298
rect -235 -307 -223 -304
rect -226 -316 -223 -307
rect -161 -313 -158 -272
rect -125 -293 -122 -271
rect 120 -290 123 -236
rect 216 -268 219 -97
rect 154 -271 219 -268
rect -132 -296 -122 -293
rect 120 -293 126 -290
rect -132 -313 -129 -296
rect -122 -313 -120 -312
rect -168 -316 -154 -313
rect -132 -316 -119 -313
rect 67 -315 81 -313
rect 123 -315 126 -293
rect 67 -316 91 -315
rect -226 -319 -214 -316
rect 78 -318 91 -316
rect 115 -318 126 -315
rect -123 -320 -121 -319
rect -244 -323 -241 -321
rect -170 -323 -120 -320
rect -244 -342 -241 -328
rect -175 -335 -172 -330
rect -176 -342 -172 -341
rect -300 -345 -172 -342
rect 20 -343 23 -331
rect 95 -343 98 -327
rect -204 -356 -201 -345
rect 20 -346 98 -343
rect 154 -346 157 -271
rect 120 -349 157 -346
rect -204 -359 -174 -356
rect -177 -403 -174 -359
rect 120 -378 123 -349
rect 37 -381 123 -378
rect -46 -403 -43 -386
rect 37 -397 40 -381
rect -177 -406 -43 -403
rect -46 -408 -43 -406
rect -1 -400 40 -397
rect -1 -408 2 -400
rect -46 -411 2 -408
<< m2contact >>
rect -162 271 -157 276
rect -321 210 -316 215
rect -158 217 -153 222
rect -321 163 -316 168
rect -236 165 -231 170
rect -256 155 -251 160
rect 99 193 104 198
rect -141 62 -136 67
rect -170 9 -165 14
rect 107 25 112 30
rect -301 -61 -296 -56
rect -162 -49 -157 -44
rect 228 85 233 90
rect 292 1 297 6
rect -129 -69 -124 -64
rect -301 -105 -296 -100
rect -296 -154 -291 -149
rect -142 -101 -136 -96
rect 98 -115 103 -110
rect -180 -148 -175 -143
rect -231 -171 -226 -166
rect -296 -198 -291 -193
rect -153 -235 -147 -230
rect -245 -283 -240 -278
rect 95 -295 100 -290
rect -245 -328 -240 -323
<< metal2 >>
rect -157 271 -46 275
rect -161 237 -156 240
rect -50 239 -46 271
rect -153 218 -49 222
rect -382 211 -321 215
rect -382 90 -378 211
rect 3 194 99 197
rect 3 182 6 194
rect -321 168 -318 169
rect -321 113 -318 163
rect -251 155 -250 160
rect -321 110 -280 113
rect -382 86 -298 90
rect -302 -56 -298 86
rect -302 -57 -301 -56
rect -350 -61 -301 -57
rect -350 -133 -346 -61
rect -283 -100 -280 110
rect -253 -40 -250 155
rect -302 -103 -301 -100
rect -296 -103 -280 -100
rect -269 -43 -250 -40
rect -292 -111 -289 -103
rect -292 -114 -278 -111
rect -350 -137 -291 -133
rect -295 -147 -291 -137
rect -337 -149 -291 -147
rect -337 -151 -296 -149
rect -337 -259 -333 -151
rect -281 -193 -278 -114
rect -291 -196 -278 -193
rect -283 -232 -280 -196
rect -269 -212 -266 -43
rect -236 -66 -233 165
rect -156 135 -153 138
rect 228 99 240 103
rect 228 90 232 99
rect -136 63 -49 67
rect 107 44 125 48
rect 107 37 111 44
rect 1 34 111 37
rect 121 36 125 44
rect 228 36 232 85
rect -120 20 -105 24
rect 1 22 4 34
rect 107 30 110 34
rect 121 32 253 36
rect 249 25 253 32
rect 249 21 296 25
rect -120 19 -112 20
rect -120 15 -116 19
rect -166 14 -116 15
rect -165 11 -116 14
rect 292 6 296 21
rect -166 -49 -162 -45
rect -236 -69 -129 -66
rect -142 -96 -49 -92
rect 87 -108 101 -105
rect 87 -109 90 -108
rect 3 -112 90 -109
rect 98 -110 101 -108
rect -142 -134 -137 -132
rect -116 -138 -110 -137
rect -119 -142 -110 -138
rect 3 -139 6 -112
rect -176 -143 -146 -142
rect -131 -143 -115 -142
rect -175 -146 -115 -143
rect -144 -147 -132 -146
rect -231 -212 -226 -171
rect -165 -192 -162 -190
rect -269 -215 -225 -212
rect -231 -230 -226 -215
rect -283 -235 -253 -232
rect -231 -235 -153 -230
rect -337 -263 -263 -259
rect -267 -274 -263 -263
rect -256 -263 -253 -235
rect -256 -266 -228 -263
rect -267 -278 -241 -274
rect -231 -323 -228 -266
rect 77 -287 98 -284
rect 10 -289 33 -288
rect 77 -289 80 -287
rect 6 -291 80 -289
rect 6 -292 14 -291
rect 25 -292 80 -291
rect 95 -290 98 -287
rect -171 -302 -110 -298
rect 6 -299 9 -292
rect -240 -326 -228 -323
rect -176 -342 -173 -341
<< m123contact >>
rect -156 236 -151 241
rect -156 130 -151 135
rect -141 24 -136 29
rect -171 -50 -166 -45
rect -142 -139 -137 -134
rect -165 -197 -160 -192
rect -176 -341 -170 -335
<< metal3 >>
rect -151 236 -62 239
rect -102 134 -99 141
rect -65 138 -62 236
rect -151 131 -99 134
rect -127 28 -40 31
rect -127 27 -124 28
rect -136 24 -124 27
rect -169 -51 -166 -50
rect -100 -51 -97 -19
rect -169 -54 -97 -51
rect -169 -55 -166 -54
rect -137 -138 -40 -134
rect -93 -193 -89 -180
rect -160 -197 -89 -193
rect -170 -339 -131 -336
rect -170 -340 -108 -339
rect -176 -342 -173 -341
rect -135 -343 -108 -340
use not  not_12
timestamp 1701035029
transform -1 0 -249 0 1 -305
box -14 -16 22 23
use not  not_8
timestamp 1701035029
transform -1 0 -140 0 1 -269
box -14 -16 22 23
use 2nand  2nand_0
timestamp 1700774385
transform -1 0 -204 0 1 -336
box -39 -3 10 38
use xor  xor_3
timestamp 1701032306
transform 1 0 -52 0 1 -286
box -69 -105 120 45
use not  not_3
timestamp 1701035029
transform 1 0 103 0 1 -316
box -14 -16 22 23
use not  not_7
timestamp 1701035029
transform -1 0 -147 0 1 -120
box -14 -16 22 23
use 3nand  3nand_0
timestamp 1700939411
transform -1 0 -181 0 1 -173
box -25 -15 34 29
use xor  xor_2
timestamp 1701032306
transform 1 0 -54 0 1 -126
box -69 -105 120 45
use not  not_2
timestamp 1701035029
transform 1 0 107 0 1 -136
box -14 -16 22 23
use not  not_5
timestamp 1701035029
transform -1 0 -146 0 1 43
box -14 -16 22 23
use 4nand  4nand_0
timestamp 1701275880
transform -1 0 -149 0 1 42
box 2 -84 80 -29
use xor  xor_1
timestamp 1701032306
transform 1 0 -54 0 1 35
box -69 -105 120 45
use not  not_1
timestamp 1701035029
transform 1 0 115 0 1 4
box -14 -16 22 23
use 5nand  5nand_0
timestamp 1701034208
transform -1 0 -193 0 1 184
box -48 -46 101 37
use xor  xor_0
timestamp 1701032306
transform 1 0 -54 0 1 195
box -69 -105 120 45
use not  not_0
timestamp 1701035029
transform 1 0 108 0 1 173
box -14 -16 22 23
use not  not_4
timestamp 1701035029
transform -1 0 -167 0 1 253
box -14 -16 22 23
use nand2  nand2_0
timestamp 1698945652
transform 1 0 248 0 1 92
box -18 -25 24 20
use not  not_11
timestamp 1701035029
transform -1 0 -300 0 1 -177
box -14 -16 22 23
use not  not_10
timestamp 1701035029
transform -1 0 -305 0 1 -84
box -14 -16 22 23
use not  not_9
timestamp 1701035029
transform -1 0 -326 0 1 184
box -14 -16 22 23
use not  not_6
timestamp 1701035029
transform 1 0 301 0 1 -37
box -14 -16 22 23
use 4nand  4nand_1
timestamp 1701275880
transform 1 0 191 0 1 34
box 2 -84 80 -29
use 4_or  4_or_0
timestamp 1699292645
transform -1 0 -377 0 1 -1
box -74 -41 134 47
<< labels >>
rlabel metal1 -517 4 -516 4 3 a_gr
rlabel metal1 327 -38 328 -38 7 equal
rlabel metal1 -127 -322 -127 -322 1 a3
rlabel metal1 -126 -315 -126 -315 1 b3
rlabel metal1 -128 -161 -128 -161 1 a2
rlabel metal1 -125 -1 -125 -1 1 a1
rlabel metal1 -127 7 -127 7 1 b1
rlabel metal1 -126 160 -126 160 1 a0
rlabel metal1 -123 168 -123 168 1 b0
rlabel metal1 51 -380 51 -380 1 gnd!
rlabel m2contact 295 3 295 3 1 vdd!
rlabel metal1 276 86 276 86 1 b_gr
rlabel metal1 -127 -154 -127 -154 1 b2
<< end >>
